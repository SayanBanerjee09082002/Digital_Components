module THIRTY_TWO_TO_FIVE_MULTIPLEXER(op, ip, s);
    input [31:0] ip;
    input [4:0] s;
    output op;
    
    assign op = (s == 5'b00000) ? ip[0] :
                (s == 5'b00001) ? ip[1] :
                (s == 5'b00010) ? ip[2] :
                (s == 5'b00011) ? ip[3] :
                (s == 5'b00100) ? ip[4] :
                (s == 5'b00101) ? ip[5] :
                (s == 5'b00110) ? ip[6] :
                (s == 5'b00111) ? ip[7] :
                (s == 5'b01000) ? ip[8] :
                (s == 5'b01001) ? ip[9] :
                (s == 5'b01010) ? ip[10] :
                (s == 5'b01011) ? ip[11] :
                (s == 5'b01100) ? ip[12] :
                (s == 5'b01101) ? ip[13] :
                (s == 5'b01110) ? ip[14] :
                (s == 5'b01111) ? ip[15] :
                (s == 5'b10000) ? ip[16] :
                (s == 5'b10001) ? ip[17] :
                (s == 5'b10010) ? ip[18] :
                (s == 5'b10011) ? ip[19] :
                (s == 5'b10100) ? ip[20] :
                (s == 5'b10101) ? ip[21] :
                (s == 5'b10110) ? ip[22] :
                (s == 5'b10111) ? ip[23] :
                (s == 5'b11000) ? ip[24] :
                (s == 5'b11001) ? ip[25] :
                (s == 5'b11010) ? ip[26] :
                (s == 5'b11011) ? ip[27] :
                (s == 5'b11100) ? ip[28] :
                (s == 5'b11101) ? ip[29] :
                (s == 5'b11110) ? ip[30] :
                ip[31];
endmodule
